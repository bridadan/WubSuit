// Actel Corporation Proprietary and Confidential
//  Copyright 2008 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
//  Revision Information:
// Jun09    Revision 4.1
// Aug10    Revision 4.2
// SVN Revision Information:
// SVN $Revision: 8508 $
// SVN $Date: 2009-06-15 16:49:49 -0700 (Mon, 15 Jun 2009) $
`timescale 1ns/1ns
module
wubsuit_base_CoreUARTapb_1_Tx_async
(
CUARTII
,
CUARTll
,
CUARTlI
,
CUARTO0I
,
CUARTI0I
,
CUARTl0I
,
CUARTOO1
,
CUARTIO1
,
CUARTlO1
,
CUARTOI1
,
CUARTII1
,
CUARTlI1
,
CUARTOl1
,
CUARTOll
)
;
parameter
TX_FIFO
=
0
;
input
CUARTII
;
input
CUARTll
;
input
CUARTlI
;
input
CUARTO0I
;
input
[
7
:
0
]
CUARTI0I
;
input
[
7
:
0
]
CUARTl0I
;
input
CUARTOO1
;
input
CUARTIO1
;
input
CUARTlO1
;
input
CUARTOI1
;
input
CUARTII1
;
output
CUARTlI1
;
wire
CUARTlI1
;
output
CUARTOl1
;
output
CUARTOll
;
reg
CUARTOl1
;
parameter
CUARTlIll
=
0
;
parameter
CUARTOlll
=
1
;
parameter
CUARTIlll
=
2
;
parameter
CUARTllll
=
3
;
parameter
CUARTO0ll
=
4
;
parameter
CUARTI0ll
=
5
;
parameter
CUARTl0ll
=
6
;
integer
CUARTO1ll
;
reg
CUARTI1ll
;
reg
[
7
:
0
]
CUARTl1ll
;
reg
[
3
:
0
]
CUARTOO0l
;
reg
CUARTIO0l
;
wire
CUARTOll
;
reg
CUARTlO0l
;
always
@
(
posedge
CUARTII
or
negedge
CUARTlI
)
begin
:
CUARTOI0l
if
(
!
CUARTlI
)
begin
CUARTI1ll
<=
1
'b
1
;
end
else
begin
if
(
TX_FIFO
==
1
'b
0
)
begin
if
(
CUARTll
)
begin
if
(
CUARTO1ll
==
CUARTIlll
)
begin
CUARTI1ll
<=
1
'b
1
;
end
end
if
(
CUARTO0I
)
begin
CUARTI1ll
<=
1
'b
0
;
end
end
else
begin
CUARTI1ll
<=
!
CUARTIO1
;
end
end
end
always
@
(
posedge
CUARTII
or
negedge
CUARTlI
)
begin
:
CUARTII0l
if
(
!
CUARTlI
)
begin
CUARTO1ll
<=
CUARTlIll
;
CUARTl1ll
<=
8
'b
0
;
CUARTlO0l
<=
1
'b
1
;
end
else
begin
if
(
CUARTll
||
(
CUARTO1ll
==
CUARTlIll
)
||
(
CUARTO1ll
==
CUARTl0ll
)
||
(
CUARTO1ll
==
CUARTOlll
)
)
begin
CUARTlO0l
<=
1
'b
1
;
case
(
CUARTO1ll
)
CUARTlIll
:
begin
if
(
TX_FIFO
==
1
'b
0
)
begin
if
(
!
CUARTI1ll
)
begin
CUARTO1ll
<=
CUARTOlll
;
end
else
begin
CUARTO1ll
<=
CUARTlIll
;
end
end
else
begin
if
(
CUARTOO1
==
1
'b
0
)
begin
CUARTlO0l
<=
1
'b
0
;
CUARTO1ll
<=
CUARTl0ll
;
end
else
begin
CUARTO1ll
<=
CUARTlIll
;
CUARTlO0l
<=
1
'b
1
;
end
end
end
CUARTOlll
:
begin
CUARTO1ll
<=
CUARTIlll
;
end
CUARTIlll
:
begin
CUARTO1ll
<=
CUARTllll
;
if
(
TX_FIFO
==
1
'b
0
)
begin
CUARTl1ll
<=
CUARTI0I
;
end
else
begin
CUARTl1ll
<=
CUARTl0I
;
end
end
CUARTllll
:
begin
if
(
CUARTlO1
)
begin
if
(
CUARTOO0l
==
4
'b
0111
)
begin
if
(
CUARTOI1
)
begin
CUARTO1ll
<=
CUARTO0ll
;
end
else
begin
CUARTO1ll
<=
CUARTI0ll
;
end
end
else
begin
CUARTO1ll
<=
CUARTllll
;
end
end
else
begin
if
(
CUARTOO0l
==
4
'b
0110
)
begin
if
(
CUARTOI1
)
begin
CUARTO1ll
<=
CUARTO0ll
;
end
else
begin
CUARTO1ll
<=
CUARTI0ll
;
end
end
else
begin
CUARTO1ll
<=
CUARTllll
;
end
end
end
CUARTO0ll
:
begin
CUARTO1ll
<=
CUARTI0ll
;
end
CUARTI0ll
:
begin
CUARTO1ll
<=
CUARTlIll
;
end
CUARTl0ll
:
begin
CUARTO1ll
<=
CUARTOlll
;
end
default
:
begin
CUARTO1ll
<=
CUARTlIll
;
end
endcase
end
end
end
assign
CUARTOll
=
CUARTlO0l
;
always
@
(
posedge
CUARTII
or
negedge
CUARTlI
)
begin
:
CUARTlI0l
if
(
!
CUARTlI
)
begin
CUARTOO0l
<=
4
'b
0000
;
end
else
begin
if
(
CUARTll
)
begin
if
(
CUARTO1ll
!=
CUARTllll
)
begin
CUARTOO0l
<=
4
'b
0000
;
end
else
begin
CUARTOO0l
<=
CUARTOO0l
+
1
'b
1
;
end
end
end
end
always
@
(
posedge
CUARTII
or
negedge
CUARTlI
)
begin
:
CUARTOl0l
if
(
!
CUARTlI
)
begin
CUARTOl1
<=
1
'b
1
;
end
else
begin
if
(
CUARTll
||
(
CUARTO1ll
==
CUARTlIll
)
||
(
CUARTO1ll
==
CUARTl0ll
)
||
(
CUARTO1ll
==
CUARTOlll
)
)
begin
case
(
CUARTO1ll
)
CUARTlIll
:
begin
CUARTOl1
<=
1
'b
1
;
end
CUARTOlll
:
begin
CUARTOl1
<=
1
'b
1
;
end
CUARTIlll
:
begin
CUARTOl1
<=
1
'b
0
;
end
CUARTllll
:
begin
CUARTOl1
<=
CUARTl1ll
[
CUARTOO0l
]
;
end
CUARTO0ll
:
begin
CUARTOl1
<=
CUARTII1
^
CUARTIO0l
;
end
CUARTI0ll
:
begin
CUARTOl1
<=
1
'b
1
;
end
default
:
begin
CUARTOl1
<=
1
'b
1
;
end
endcase
end
end
end
always
@
(
posedge
CUARTII
or
negedge
CUARTlI
)
begin
:
CUARTIl0l
if
(
!
CUARTlI
)
begin
CUARTIO0l
<=
1
'b
0
;
end
else
begin
if
(
CUARTll
&
CUARTOI1
)
begin
if
(
CUARTO1ll
==
CUARTllll
)
begin
CUARTIO0l
<=
CUARTIO0l
^
CUARTl1ll
[
CUARTOO0l
]
;
end
else
begin
CUARTIO0l
<=
CUARTIO0l
;
end
end
if
(
CUARTO1ll
==
CUARTI0ll
)
begin
CUARTIO0l
<=
1
'b
0
;
end
end
end
assign
CUARTlI1
=
CUARTI1ll
;
endmodule
